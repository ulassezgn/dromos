package control_pkg;
    typedef enum logic [2:0] {
        R_TYPE;
        I_TYPE;
        S_TYPE;
        B_TYPE;
        U_TYPE;
        J_TYPE;
    } instr_type_e;

endpackage